package packet_pkg;
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/packet_data.sv"
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/component_base.sv"
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/sequencer.sv"
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/driver.sv"
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/monitor.sv"
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/agent.sv"
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/packet_vc.sv"
	//`include "/data.cc/data/a/home/cc/students/enginer/yazanatamna/project_leen_yazan/checker.sv"
endpackage