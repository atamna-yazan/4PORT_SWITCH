module top_test;
import packet_pkg::*;
switch_test test_h();   
endmodule
