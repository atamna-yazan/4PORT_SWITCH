class packet;
	logic [3:0] source;
	logic [3:0] target;
	logic [7:0] data;

	function new(string n="pkt");
	endfunction
  endclass